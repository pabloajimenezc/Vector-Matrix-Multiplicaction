magic
tech sky130A
timestamp 1702662493
<< nwell >>
rect 2600 -500 5200 2400
<< nmos >>
rect 3900 -1800 4000 -1300
<< pmos >>
rect 3900 -100 4000 1400
<< ndiff >>
rect 3200 -1400 3900 -1300
rect 3200 -1700 3300 -1400
rect 3500 -1700 3900 -1400
rect 3200 -1800 3900 -1700
rect 4000 -1400 4700 -1300
rect 4000 -1700 4400 -1400
rect 4600 -1700 4700 -1400
rect 4000 -1800 4700 -1700
<< pdiff >>
rect 3200 1200 3900 1400
rect 3200 900 3300 1200
rect 3500 900 3900 1200
rect 3200 -100 3900 900
rect 4000 1200 4700 1400
rect 4000 900 4400 1200
rect 4600 900 4700 1200
rect 4000 -100 4700 900
<< ndiffc >>
rect 3300 -1700 3500 -1400
rect 4400 -1700 4600 -1400
<< pdiffc >>
rect 3300 900 3500 1200
rect 4400 900 4600 1200
<< poly >>
rect 3900 1400 4000 1500
rect 3900 -700 4000 -100
rect 3300 -800 4000 -700
rect 3300 -1000 3400 -800
rect 3800 -1000 4000 -800
rect 3300 -1100 4000 -1000
rect 3900 -1300 4000 -1100
rect 3900 -1900 4000 -1800
<< polycont >>
rect 3400 -1000 3800 -800
<< locali >>
rect 2900 1700 4900 2000
rect 3200 1200 3500 1700
rect 3200 900 3300 1200
rect 3200 -100 3500 900
rect 4400 1200 4700 1400
rect 4600 900 4700 1200
rect 3300 -800 3900 -700
rect 3300 -1000 3400 -800
rect 3800 -1000 3900 -800
rect 3300 -1100 3900 -1000
rect 3200 -1400 3500 -1300
rect 3200 -1700 3300 -1400
rect 3200 -2200 3500 -1700
rect 4400 -1400 4700 900
rect 4600 -1700 4700 -1400
rect 4400 -1800 4700 -1700
rect 2900 -2500 4900 -2200
<< metal1 >>
rect 2700 1400 5100 2300
rect 2700 -2800 5100 -1900
<< end >>
